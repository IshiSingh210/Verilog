module MUX_16(S3,S2,S1,S0,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,Y);
  input S3,S2,S1,S0,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15;
  output Y;
  assign Y=(~S3&~S2&~S1&~S0&I0)|(~S3&~S2&~S1&S0&I1)|(~S3&~S2&S1&~S0&I2)|(~S3&~S2&S1&S0&I3)|(~S3&S2&~S1&~S0&I4)
  |(~S3&S2&~S1&S0&I5)|(~S3&S2&S1&~S0&I6)|(~S3&S2&S1&S0&I7)|(S3&~S2&~S1&~S0&I8)|(S3&~S2&~S1&S0&I9)
  |(S3&~S2&S1&~S0&I10)|(S3&~S2&S1&S0&I11)|(S3&S2&~S1&~S0&I12)|(S3&S2&~S1&S0&I13)|(S3&S2&S1&~S0&I4)|(S3&S2&S1&S0&I15);
endmodule

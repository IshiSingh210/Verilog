module BCDripple(clr,clk,dir, tc, q);
input clr,clk,dir;
output reg tc;
output reg[3:0] q;
always@(posedge clk,posedge clr)
begin
  if(clr==1)
    q=4'd0;
  else
    begin
      if (dir==1)
        q=q+1;
      else if(dir==0)
        q=q-1;
      if(dir==1 & q==4'd10) 
      begin
        q=4'd0;
        tc=1'b1;
      end
      else if(dir==0 & q==4'd15)
      begin
        q=1'd9;
        tc=1'b1;
      end
      else 
        tc=1'b0;  
    end
end 
endmodule